module io();

endmodule